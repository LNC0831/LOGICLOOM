module ALU (clk, rst, cmd, input1, input2, \output );
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] cmd;
  input  wire [7:0] input1;
  input  wire [7:0] input2;
  output  wire [7:0] \output ;

  TC_Or # (.UUID(64'd1029278905383820776 ^ UUID), .BIT_WIDTH(64'd8)) Or8_0 (.in0(wire_20), .in1(wire_31), .out(wire_16));
  TC_Not # (.UUID(64'd1855087917867058098 ^ UUID), .BIT_WIDTH(64'd8)) Not8_1 (.in(wire_18), .out(wire_20));
  TC_Not # (.UUID(64'd1120555654468192161 ^ UUID), .BIT_WIDTH(64'd8)) Not8_2 (.in(wire_14), .out(wire_31));
  TC_Or # (.UUID(64'd4087604044960771246 ^ UUID), .BIT_WIDTH(64'd8)) Or8_3 (.in0(wire_34), .in1(wire_22), .out(wire_21));
  TC_Not # (.UUID(64'd1605617921455847448 ^ UUID), .BIT_WIDTH(64'd8)) Not8_4 (.in(wire_21), .out(wire_30));
  TC_Or # (.UUID(64'd2585052386329273930 ^ UUID), .BIT_WIDTH(64'd8)) Or8_5 (.in0(wire_37), .in1(wire_17), .out(wire_36));
  TC_Not # (.UUID(64'd3425828984370853204 ^ UUID), .BIT_WIDTH(64'd8)) Not8_6 (.in(wire_36), .out(wire_25));
  TC_Not # (.UUID(64'd673144019471828146 ^ UUID), .BIT_WIDTH(64'd8)) Not8_7 (.in(wire_26), .out(wire_37));
  TC_Not # (.UUID(64'd3365265557724810005 ^ UUID), .BIT_WIDTH(64'd8)) Not8_8 (.in(wire_10), .out(wire_17));
  TC_Or # (.UUID(64'd3577820485719657908 ^ UUID), .BIT_WIDTH(64'd8)) Or8_9 (.in0(wire_19), .in1(wire_28), .out(wire_23));
  TC_Splitter8 # (.UUID(64'd2795288827045885747 ^ UUID)) Splitter8_10 (.in(wire_35), .out0(wire_32), .out1(wire_24), .out2(wire_29), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd4468983803232351222 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_0), .in(wire_4), .out(wire_18));
  TC_Switch # (.UUID(64'd395591505664693870 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_0), .in(wire_9), .out(wire_14));
  TC_Switch # (.UUID(64'd1601402203432394550 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_3), .in(wire_4), .out(wire_34));
  TC_Switch # (.UUID(64'd970195613402418433 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_14 (.en(wire_3), .in(wire_9), .out(wire_22));
  TC_Switch # (.UUID(64'd1974079933648512979 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_8), .in(wire_4), .out(wire_26));
  TC_Switch # (.UUID(64'd2113715048216053677 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_8), .in(wire_9), .out(wire_10));
  TC_Switch # (.UUID(64'd1417111000291069272 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_7), .in(wire_4), .out(wire_19));
  TC_Switch # (.UUID(64'd2620733236984203592 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_7), .in(wire_9), .out(wire_28));
  TC_Decoder3 # (.UUID(64'd3431927245054413885 ^ UUID)) Decoder3_19 (.dis(1'd0), .sel0(wire_32), .sel1(wire_24), .sel2(wire_29), .out0(wire_7), .out1(wire_0), .out2(wire_3), .out3(wire_8), .out4(wire_6), .out5(wire_5), .out6(), .out7());
  TC_Switch # (.UUID(64'd888147644563154846 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_20 (.en(wire_7), .in(wire_23), .out(wire_2_1));
  TC_Switch # (.UUID(64'd2228716300505859704 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_21 (.en(wire_0), .in(wire_16), .out(wire_2_0));
  TC_Switch # (.UUID(64'd1607598335967245297 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_22 (.en(wire_3), .in(wire_30), .out(wire_2_2));
  TC_Switch # (.UUID(64'd299260152923995108 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_23 (.en(wire_8), .in(wire_25), .out(wire_2_3));
  TC_Add # (.UUID(64'd169074278508500186 ^ UUID), .BIT_WIDTH(64'd8)) Add8_24 (.in0(wire_1), .in1(wire_11), .ci(1'd0), .out(wire_15), .co());
  TC_Add # (.UUID(64'd2574134166858126510 ^ UUID), .BIT_WIDTH(64'd8)) Add8_25 (.in0(wire_27), .in1(wire_12), .ci(1'd0), .out(wire_33), .co());
  TC_Switch # (.UUID(64'd629117182162894566 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_26 (.en(wire_6), .in(wire_4), .out(wire_1));
  TC_Switch # (.UUID(64'd4347130703739876119 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_27 (.en(wire_6), .in(wire_9), .out(wire_11));
  TC_Switch # (.UUID(64'd2731706839471440459 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_28 (.en(wire_6), .in(wire_15), .out(wire_2_4));
  TC_Neg # (.UUID(64'd1635506308924341396 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_29 (.in(wire_13), .out(wire_12));
  TC_Switch # (.UUID(64'd2718341691260391934 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_30 (.en(wire_5), .in(wire_4), .out(wire_27));
  TC_Switch # (.UUID(64'd1850747926098071791 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_31 (.en(wire_5), .in(wire_9), .out(wire_13));
  TC_Switch # (.UUID(64'd1099209684752076663 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_32 (.en(wire_5), .in(wire_33), .out(wire_2_5));

  wire [0:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_2_0;
  wire [7:0] wire_2_1;
  wire [7:0] wire_2_2;
  wire [7:0] wire_2_3;
  wire [7:0] wire_2_4;
  wire [7:0] wire_2_5;
  assign wire_2 = wire_2_0|wire_2_1|wire_2_2|wire_2_3|wire_2_4|wire_2_5;
  assign \output  = wire_2;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  assign wire_4 = input1;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [7:0] wire_9;
  assign wire_9 = input2;
  wire [7:0] wire_10;
  wire [7:0] wire_11;
  wire [7:0] wire_12;
  wire [7:0] wire_13;
  wire [7:0] wire_14;
  wire [7:0] wire_15;
  wire [7:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_18;
  wire [7:0] wire_19;
  wire [7:0] wire_20;
  wire [7:0] wire_21;
  wire [7:0] wire_22;
  wire [7:0] wire_23;
  wire [0:0] wire_24;
  wire [7:0] wire_25;
  wire [7:0] wire_26;
  wire [7:0] wire_27;
  wire [7:0] wire_28;
  wire [0:0] wire_29;
  wire [7:0] wire_30;
  wire [7:0] wire_31;
  wire [0:0] wire_32;
  wire [7:0] wire_33;
  wire [7:0] wire_34;
  wire [7:0] wire_35;
  assign wire_35 = cmd;
  wire [7:0] wire_36;
  wire [7:0] wire_37;

endmodule
