module CPU (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_Splitter8 # (.UUID(64'd1740909036157118627 ^ UUID)) Splitter8_0 (.in(wire_6), .out0(wire_16), .out1(wire_4), .out2(wire_34), .out3(wire_11), .out4(wire_17), .out5(wire_19), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd3285532197686644414 ^ UUID)) Decoder3_1 (.dis(wire_31), .sel0(wire_16), .sel1(wire_4), .sel2(wire_34), .out0(wire_21), .out1(wire_36), .out2(wire_26), .out3(wire_28), .out4(wire_10), .out5(wire_22), .out6(wire_9), .out7());
  TC_Decoder3 # (.UUID(64'd2068417560946943622 ^ UUID)) Decoder3_2 (.dis(wire_31), .sel0(wire_11), .sel1(wire_17), .sel2(wire_19), .out0(wire_18), .out1(wire_29), .out2(wire_8), .out3(wire_20), .out4(wire_32), .out5(wire_27), .out6(wire_3), .out7());
  TC_Switch # (.UUID(64'd325150327384652478 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_3 (.en(wire_5), .in(wire_30), .out(wire_2_8));
  TC_Mux # (.UUID(64'd723863209402855404 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_4 (.sel(wire_5), .in0({{7{1'b0}}, wire_28 }), .in1({{7{1'b0}}, wire_5 }), .out(wire_37));
  TC_Counter # (.UUID(64'd2647770476147775263 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_5 (.clk(clk), .rst(rst), .save(wire_1), .in(wire_12), .out(wire_13));
  TC_Mux # (.UUID(64'd4158782181600309462 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_6 (.sel(wire_15), .in0({{7{1'b0}}, wire_21 }), .in1({{7{1'b0}}, wire_15 }), .out(wire_7));
  TC_Switch # (.UUID(64'd3888359016934678901 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_15), .in(wire_6), .out(wire_2_0));
  TC_Not # (.UUID(64'd3155310201563455113 ^ UUID), .BIT_WIDTH(64'd1)) Not_8 (.in(wire_0), .out(wire_31));
  TC_Switch # (.UUID(64'd347437319060339452 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_9 (.en(wire_23), .in(wire_6), .out(wire_35));
  TC_Program8_1 # (.UUID(64'd857501675760812171 ^ UUID), .DEFAULT_FILE_NAME("Program8_1_BE6753B1A06808B.w8.bin"), .ARG_SIG("Program8_1_BE6753B1A06808B=%s")) Program8_1_10 (.clk(clk), .rst(rst), .address(wire_13), .out(wire_6));
  TC_Switch # (.UUID(64'd1502156430737279918 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_3), .in(wire_24), .out(wire_2_2));
  TC_Constant # (.UUID(64'd1643049279126162415 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5)) Constant8_12 (.out(wire_24));
  TC_SegmentDisplay # (.UUID(64'd4193781903170062915 ^ UUID)) SegmentDisplay_13 (.clk(clk), .rst(rst), .enable(wire_9), .value(wire_2));
  DEC # (.UUID(64'd561234129375555341 ^ UUID)) DEC_14 (.clk(clk), .rst(rst), .opcode(wire_6), .imme(wire_15), .condition(wire_23), .cal(wire_5), .copy(wire_0));
  ALU # (.UUID(64'd3203376692861713137 ^ UUID)) ALU_15 (.clk(clk), .rst(rst), .cmd(wire_6), .input1(wire_25), .input2(wire_14), .\output (wire_30));
  COND # (.UUID(64'd3319144537462594360 ^ UUID)) COND_16 (.clk(clk), .rst(rst), .condition(wire_35), .\input (wire_33), .\output (wire_1));
  RegisterPlus # (.UUID(64'd2013824320296903733 ^ UUID)) RegisterPlus_17 (.clk(clk), .rst(rst), .rd_en(wire_18), .\input (wire_2), .wr_en(wire_7[0:0]), .output_always(wire_12), .Output(wire_2_7));
  RegisterPlus # (.UUID(64'd4393917700000120423 ^ UUID)) RegisterPlus_18 (.clk(clk), .rst(rst), .rd_en(wire_29), .\input (wire_2), .wr_en(wire_36), .output_always(wire_25), .Output(wire_2_6));
  RegisterPlus # (.UUID(64'd898038243217137729 ^ UUID)) RegisterPlus_19 (.clk(clk), .rst(rst), .rd_en(wire_8), .\input (wire_2), .wr_en(wire_26), .output_always(wire_14), .Output(wire_2_5));
  RegisterPlus # (.UUID(64'd2922266585936576169 ^ UUID)) RegisterPlus_20 (.clk(clk), .rst(rst), .rd_en(wire_20), .\input (wire_2), .wr_en(wire_37[0:0]), .output_always(wire_33), .Output(wire_2_4));
  RegisterPlus # (.UUID(64'd2122138527428093258 ^ UUID)) RegisterPlus_21 (.clk(clk), .rst(rst), .rd_en(wire_32), .\input (wire_2), .wr_en(wire_10), .output_always(), .Output(wire_2_3));
  RegisterPlus # (.UUID(64'd4446153895860665334 ^ UUID)) RegisterPlus_22 (.clk(clk), .rst(rst), .rd_en(wire_27), .\input (wire_2), .wr_en(wire_22), .output_always(), .Output(wire_2_1));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_2_0;
  wire [7:0] wire_2_1;
  wire [7:0] wire_2_2;
  wire [7:0] wire_2_3;
  wire [7:0] wire_2_4;
  wire [7:0] wire_2_5;
  wire [7:0] wire_2_6;
  wire [7:0] wire_2_7;
  wire [7:0] wire_2_8;
  assign wire_2 = wire_2_0|wire_2_1|wire_2_2|wire_2_3|wire_2_4|wire_2_5|wire_2_6|wire_2_7|wire_2_8;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [7:0] wire_6;
  wire [7:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [7:0] wire_12;
  wire [7:0] wire_13;
  wire [7:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [7:0] wire_24;
  wire [7:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [7:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [7:0] wire_33;
  wire [0:0] wire_34;
  wire [7:0] wire_35;
  wire [0:0] wire_36;
  wire [7:0] wire_37;

endmodule
